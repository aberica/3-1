// memwb_reg.v
// This module is the MEM/WB pipeline register.


module memwb_reg #(
  parameter DATA_WIDTH = 32
)(
  // TODO: Add flush or stall signal if it is needed

  //////////////////////////////////////
  // Inputs
  //////////////////////////////////////
  input clk,

  input [DATA_WIDTH-1:0] mem_pc_plus_4,

  // wb control
  input [1:0] mem_jump,
  input mem_memtoreg,
  input mem_regwrite,
  
  input [DATA_WIDTH-1:0] mem_readdata,
  input [DATA_WIDTH-1:0] mem_alu_result,
  input [4:0] mem_rd,
  
  //////////////////////////////////////
  // Outputs
  //////////////////////////////////////
  output [DATA_WIDTH-1:0] wb_pc_plus_4,

  // wb control
  output [1:0] wb_jump,
  output wb_memtoreg,
  output wb_regwrite,
  
  output [DATA_WIDTH-1:0] wb_readdata,
  output [DATA_WIDTH-1:0] wb_alu_result,
  output [4:0] wb_rd
);

// TODO: Implement MEM/WB pipeline register module
  // Reg
  reg [DATA_WIDTH-1:0] wb_pc_plus_4_reg;

  // wb control
  reg [1:0] wb_jump_reg;
  reg wb_memtoreg_reg;
  reg wb_regwrite_reg;
  
  reg [DATA_WIDTH-1:0] wb_readdata_reg;
  reg [DATA_WIDTH-1:0] wb_alu_result_reg;
  reg [4:0] wb_rd_reg;


  // Assign
  assign wb_pc_plus_4 = wb_pc_plus_4_reg;

  // wb control
  assign wb_jump = wb_jump_reg;
  assign wb_memtoreg = wb_memtoreg_reg;
  assign wb_regwrite = wb_regwrite_reg;

  assign wb_readdata = wb_readdata_reg;
  assign wb_alu_result = wb_alu_result_reg;
  assign wb_rd = wb_rd_reg;


  always @(posedge clk) begin
    wb_pc_plus_4_reg <= mem_pc_plus_4;

    // wb control
    wb_jump_reg <= mem_jump;
    wb_memtoreg_reg <= mem_memtoreg;
    wb_regwrite_reg <= mem_regwrite;

    wb_readdata_reg <= mem_readdata;
    wb_alu_result_reg <= mem_alu_result;
    wb_rd_reg <= mem_rd;
  end

endmodule
